library verilog;
use verilog.vl_types.all;
entity freq_divider_vlg_vec_tst is
end freq_divider_vlg_vec_tst;
